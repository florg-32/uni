//=============================================================================
// Project  : Industrial HW Verification
//
// File Name: avmm_sequencer.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2016-04-18-EP on Thu Apr 28 06:08:21 2022
//=============================================================================
// Description: Sequencer for avmm
//=============================================================================

`ifndef AVMM_SEQUENCER_SV
`define AVMM_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(avmm_tr) avmm_sequencer_t;


`endif // AVMM_SEQUENCER_SV

